module memory_system_testbench();

endmodule