module alu_testbench();

endmodule