module full_system_testbench();


endmodule