module memory_controller_testbench();


endmodule