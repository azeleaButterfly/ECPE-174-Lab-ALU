module memory_module_testbench();


endmodule